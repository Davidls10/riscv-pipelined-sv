module instruction_memory(input logic [31:0] pc,
                          output logic [31:0] instr);

    /*
    L1: lw x5, -4(x9)        I   111111111100 01001 010 00101 0000011 // stall when in the execute stage
        or x4, x5, x6        R   0000000 00110 00101 110 00100 0110011 // forwarding
        sw x6, 8(x9)         S   0000000 00110 01001 010 01000 0100011 // normal
        addi x4, x4, 2       I   000000000010 00100 000 00100 0010011 // forwarding
        sw x4, 4(x9)         S   0000000 00100 01001 010 00100 0100011 // normal
        lw x5, 4(x9)         I   000000000100 01001 010 00101 0000011 // stall
        and x4, x4, x5       R   0000000 00101 00100 111 00100 0110011 // forwarding
        beq x4, x5, L1       B   1111111 00101 00100 000 00101 1100011 // FlushD
    */

    always_comb begin
        case(pc)
            32'h0000: instr = 32'b11111111110001001010001010000011;
            32'h0004: instr = 32'b00000000011000101110001000110011;
            32'h0008: instr = 32'b00000000011001001010010000100011;
            32'h000c: instr = 32'b00000000001000100000001000010011;
            32'h0010: instr = 32'b00000000010001001010001000100011;
            32'h0014: instr = 32'b00000000010001001010001010000011;
            32'h0018: instr = 32'b00000000010100100111001000110011;
            32'h001c: instr = 32'b11111110010100100000001011100011;

            default:  instr = 32'b0;
        endcase
    end
    
endmodule
